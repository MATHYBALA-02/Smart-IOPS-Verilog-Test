module andgate(
	input a,b,
	output c);
c=a and b;
$display("the output is %d",c);
endmodule
